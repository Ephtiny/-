module vending_machine(
	input  wire 		 clk,//??
	input  wire 		 rst_n,//??
	input        [3:0] key_value,//???
	input        [3:0] flag,
	
	output reg        beep,
	output reg   [3:0] led,
	output wire   [3:0] money_flag_w,
	output wire  boot_flag_w
);

parameter MAX_NUM = 9_999_999;//??????0.2s  LED?????
parameter MAX_NUM2 = 10;//2s????0.2s

//????????4??4???
reg [1:0] led_flag; 

reg boot_flag;                   //????????????? 0??? 1???

reg [3:0] money_flag;//????????8? ???0, 0.5, 1, 1.5, 2, 2.5, 3, 3.5, ???0

reg [23:0] cnt = 0;             //???????0

reg [26:0] cnt_1 = 0;             //???????0

reg time_flag;//?????? 1:???? 0:???



//0.2s?????
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)
		cnt <= 1'b0;               //????????
	else if(cnt == MAX_NUM)          //???????????????
      cnt <= 1'b0;
	else
		cnt <= cnt + 1'b1;         
end

//2s?????
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)
		cnt_1 <= 1'b0;               //????????
	else if(time_flag == 1)begin//????
		if(cnt == MAX_NUM)begin
			if(cnt_1 <MAX_NUM2)begin
				cnt_1 <= cnt_1 + 1'b1;
			end
			else begin
				cnt_1 <= 1'b0;//cnt_1?????????
			end
		end
		else begin
			cnt_1 <= cnt_1;//??????
		end
	end
	else begin
		cnt_1 <= 1'b0;//????cnt_1??
	end
end


//????????? led_flag?????0.2s
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)
		led_flag <= 1'b0;
	else if(cnt == MAX_NUM)
		led_flag <= led_flag + 1'b1;      //?????????
	else
		led_flag <= led_flag;
end 


//?????????? key4
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)begin  
			boot_flag <= 1'b0;                 //???????
			beep <= 1'b0;//????????? 
	end
	else if(flag[3] == 1'b1 && key_value[3] == 1'b0)begin//???key4??????????????
			boot_flag <= ~boot_flag;
			beep <= ~beep;//???????????
		end
	else begin
		boot_flag <= boot_flag;//??????????????
		beep <= beep;//???????
	end
end


assign boot_flag_w = boot_flag;

//??????????
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)begin
		money_flag <= 4'd0;//???????0
	end
	else if(boot_flag)begin//????????????????
		case(money_flag)
			4'd0:begin//?????0????
				if(flag[1] == 1'b1 && key_value[1] == 1'b0)begin//????0.5
					money_flag <= 4'd1;//???????
				end
				else if(flag[2] == 1'b1 && key_value[2] == 1'b0)begin//????1
					money_flag <= 4'd2;//???????
				end
//				else if(flag[0] == 1'b1 && key_value[0] == 1'b0)begin//????
//					money_flag <= 4'd7;//???????
//					time_flag <= 1'b1;//????
//				end
				else begin//??????????
					money_flag <= money_flag;
				end
			end
			4'd1:begin//?????0.5????
				if(flag[1] == 1'b1 && key_value[1] == 1'b0)begin//????0.5
					money_flag <= 4'd2;//???????
				end
				else if(flag[2] == 1'b1 && key_value[2] == 1'b0)begin//????1
					money_flag <= 4'd3;//???????
				end
				else if(flag[0] == 1'b1 && key_value[0] == 1'b0)begin//????
				money_flag <= 4'd7;//???????
				time_flag <= 1'b1;//????
				end
				else begin//??????????
					money_flag <= money_flag;
				end
			end
			4'd2:begin//?????1????
				if(flag[1] == 1'b1 && key_value[1] == 1'b0)begin//????0.5
					money_flag <= 4'd3;//???????
				end
				else if(flag[2] == 1'b1 && key_value[2] == 1'b0)begin//????1
					money_flag <= 4'd4;//???????
				end
				else if(flag[0] == 1'b1 && key_value[0] == 1'b0)begin//????
					money_flag <= 4'd7;//???????
					time_flag <= 1'b1;//????
				end
				else begin//??????????
					money_flag <= money_flag;
				end
			end
			4'd3:begin//?????1.5????
				if(flag[1] == 1'b1 && key_value[1] == 1'b0)begin//????0.5
					money_flag <= 4'd4;//???????
				end
				else if(flag[2] == 1'b1 && key_value[2] == 1'b0)begin//????1
					money_flag <= 4'd5;//???????
					time_flag <= 1'b1;//????
				end
				else if(flag[0] == 1'b1 && key_value[0] == 1'b0)begin//????
					money_flag <= 4'd7;//???????
					time_flag <= 1'b1;//????
				end
				else begin//??????????
					money_flag <= money_flag;
				end
			end
			4'd4:begin//?????2????
				if(flag[1] == 1'b1 && key_value[1] == 1'b0)begin//????0.5
					money_flag <= 4'd5;//???????
					time_flag <= 1'b1;//????
				end
				else if(flag[2] == 1'b1 && key_value[2] == 1'b0)begin//????1
					money_flag <= 4'd6;//???????
					time_flag <= 1'b1;//????
				end
				else if(flag[0] == 1'b1 && key_value[0] == 1'b0)begin//????
					money_flag <= 4'd7;//???????
					time_flag <= 1'b1;//????
				end
				else begin//??????????
					money_flag <= money_flag;
				end
			end
			4'd5:begin//?????2.5???? ??2s
				if(cnt_1 == MAX_NUM2)begin
					money_flag <= 4'd0;//???????
					time_flag <= 1'b0;//????
				end
				else begin
					money_flag <= money_flag;
				end
			end
			4'd6:begin//?????3???? ??2s
				if(cnt_1 == MAX_NUM2)begin
					money_flag <= 4'd0;//???????
					time_flag <= 1'b0;//????
				end
				else begin
					money_flag <= money_flag;
				end
			end
			4'd7:begin//???????? ??2s
				if(cnt_1 == MAX_NUM2)begin
					money_flag <= 4'd0;//???????
					time_flag <= 1'b0;//????
				end
				else begin
					money_flag <= money_flag;
				end
			end
		endcase
	end
	else begin
		money_flag <= 4'd0;
	end
end




//led????
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)
		led <= 4'b0000;
	else if(money_flag == 4'd5)begin//2.5????????  ??
			case(led_flag)
				2'b00  :led <= 4'b1111;
				2'b01  :led <= 4'b0000;
				2'b10  :led <= 4'b1111;
				2'b11  :led <= 4'b0000;
				default:led <= 4'b1111;
			endcase
	end
	else if(money_flag == 4'd6)begin//3???????  ???
			case(led_flag)
				2'b00  :led <= 4'b1000;
				2'b01  :led <= 4'b0100;
				2'b10  :led <= 4'b0010;
				2'b11  :led <= 4'b0001;
				default:led <= 4'b1000;
			endcase
	end
	else if(money_flag == 4'd7)begin//?? ????????
			case(led_flag)
				2'b00  :led <= 4'b1000;
				2'b01  :led <= 4'b1100;
				2'b10  :led <= 4'b1110;
				2'b11  :led <= 4'b1111;
				default:led <= 4'b1000;
			endcase
	end
	else
		led <= 4'b0000;//????led??
end


assign money_flag_w = money_flag;

endmodule