module my_vending_machine(
	input	logic	      clk,
	input	logic	      rst_n,  // ???
    	input	logic	[2:0] key_value,  // ???

	output	logic	      beep,  // ??&????
    	output	logic	[3:0] money_flag  // ????
);
    
    parameter ts = 20'd3_999;  // ???????
    
    logic  [19:0] cnt = 0;  // ??????
    
    always @(posedge clk or negedge rst_n)
        begin
            if (!rst_n) begin
                cnt <= 20'd0;
                beep <= 0;
                money_flag <= 4'd0;
            end
            else
                cnt = cnt + 1;
        end
    
    always @(*)
        begin
            if (cnt == ts) begin
                case(money_flag)
                    4'd0:begin
                	money_flag = 4'd0;
                    end
                    default:begin
                	money_flag <= 4'd7;
                	cnt <= 20'd0;
                    end
                endcase
	    end
	    else begin
		money_flag = money_flag;
	    end
	end
                        
    always @(posedge clk or negedge clk)
        begin
            case(money_flag)
                4'd0:begin//?????0????
			beep <= 0;
			if(key_value[1] == 1'b0)begin//????0.5
				money_flag <= 4'd1;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[2] == 1'b0)begin//????1
				money_flag <= 4'd2;//???????
                      		cnt <= 20'd0;
			end
                  	else begin
                      		money_flag <= money_flag;
                  	end
		end
		4'd1:begin//?????0.5????
			if(key_value[1] == 1'b0)begin//????0.5
				money_flag <= 4'd2;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[2] == 1'b0)begin//????1
				money_flag <= 4'd3;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[0] == 1'b0)begin//????
				money_flag <= 4'd7;//???????
                      		cnt <= 20'd0;
			end
                  	else begin
                      		money_flag <= money_flag;
                  	end
		end
		4'd2:begin//?????1????
			if(key_value[1] == 1'b0)begin//????0.5
				money_flag <= 4'd3;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[2] == 1'b0)begin//????1
				money_flag <= 4'd4;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[0] == 1'b0)begin//????
				money_flag <= 4'd7;//???????
                      		cnt <= 20'd0;
			end
                  	else begin
                      		money_flag <= money_flag;
                  	end
		end
		4'd3:begin//?????1.5????
			if(key_value[1] == 1'b0)begin//????0.5
				money_flag <= 4'd4;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[2] == 1'b0)begin//????1
				money_flag <= 4'd5;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[0] == 1'b0)begin//????
				money_flag <= 4'd7;//???????
                      		cnt <= 20'd0;
			end
                  	else begin
                      		money_flag <= money_flag;
                  	end
		end
		4'd4:begin//?????2????
			if(key_value[1] == 1'b0)begin//????0.5
				money_flag <= 4'd5;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[2] == 1'b0)begin//????1
				money_flag <= 4'd6;//???????
                      		cnt <= 20'd0;
			end
			else if(key_value[0] == 1'b0)begin//????
				money_flag <= 4'd7;//???????
                      		cnt <= 20'd0;
			end
                  	else begin
                      	money_flag <= money_flag;
                  	end
		end
		4'd5:begin//?????2.5????
			money_flag <= 4'd0;  // ??????????
		end
		4'd6:begin//?????3????
			money_flag <= 4'd0;  // ??????????
			beep <= 1;  // ??
		end
		4'd7:begin//????????
			money_flag <=4'd0;
                	beep = 1;
		end
            endcase
        end
endmodule
