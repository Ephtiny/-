module key_debounce(
	input  wire  clk,
	input  wire  rst_n,
	input  wire  key,
	
	output reg   flag,               //??????????????0????1?????
	output reg   key_value           //????????????????
);

//??20ms?????,0.2s,1_000_000?
reg [19:0] delay_cnt;

//????key??????????????
reg key_reg;



//20ms?????
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)
		begin
			key_reg <= 1'b1;                        //???????????
			delay_cnt <= 1'b0;                      //??????0
		end
	else
		begin
			key_reg <= key; 
			if(key_reg == 1 && key == 0)            //????key?????key???????????
				delay_cnt <= 20'd1_000_000;          //????20ms
			else if(delay_cnt > 0)
				delay_cnt <= delay_cnt - 1;          //???????20ms???
			else
				delay_cnt <= 1'b0;                  
		end
end


//??????????????????
always@(posedge clk or negedge rst_n)begin
	if(!rst_n)
		begin
		   flag <= 1'b0;                               //??????????????
			key_value <= 1'b1;                          //??????1
		end
	else
		begin
			if(delay_cnt == 20'd1)                      //???1_000_000?1
				begin
					flag <= 1'b1;
					key_value <= key;                     //??20ms??key???key_value
				end
			else	
				begin
					flag <= 1'b0;
					key_value <= key_value;               //20ms?????
				end
		end
end

endmodule
